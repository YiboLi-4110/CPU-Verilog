`ifndef ALUOp_DEFS
`define ALUOp_DEFS

`define ALUOp_WIRENUM   4

`define ALUOp_ADD       4'b0000
`define ALUOp_SUB       4'b0001
`define ALUOp_ADDU      4'b0010
`define ALUOp_SUBU      4'b0011
`define ALUOp_SLT       4'b0100
`define ALUOp_SLTU      4'b0101
`define ALUOp_AND       4'b0110
`define ALUOp_OR        4'b0111
`define ALUOp_XOR       4'b1000
`define ALUOp_R         4'b1111

`endif