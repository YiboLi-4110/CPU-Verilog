`ifndef OP_CODE
`define OP_CODE

`define OP_CODE_LW 6'b100011
`define OP_CODE_SW 6'b101011
`define OP_CODE_RR 6'b000000
`define OP_CODE_ADDI 6'b001000
`define OP_CODE_ADDIU 6'b001001
`define OP_CODE_ANDI 6'b001100
`define OP_CODE_ORI 6'b001101
`define OP_CODE_XORI 6'b001110
`define OP_CODE_SLTI 6'b001010
`define OP_CODE_SLTIU 6'b001011
`define OP_CODE_BEQ 6'b000100
`define OP_CODE_BNE 6'b000101
`define OP_CODE_BLEZ 6'b000110
`define OP_CODE_BGTZ 6'b000111
`define OP_CODE_BLTZ 6'b000001
`define OP_CODE_BGEZ 6'b000001
`define OP_CODE_J 6'b000010
`define OP_CODE_JAL 6'b000011
`define OP_CODE_LUI 6'b001111

`endif 